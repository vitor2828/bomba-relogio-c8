module counter (input logic clk
                input logic reset
                output logic [5:0]q);

always_ff @(posedge clk, posedge reset)
    if (reset)
        q <= 0;
    else begin
        q <= q + 1;

endmodule