module register_senha_B (
	input logic clk,
	input logic en,
	input logic [2:0] d,
	output logic [2:0] q
);

	always_ff@(posedge clk, posedge en) begin
		if (en) begin
			q <= d;
		end
	end
		
endmodule

